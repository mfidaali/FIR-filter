//////////////////////////////////////////////////////////////////////
////                                                              ////
//// registerInterface.v                                          ////
////                                                              ////
//// This file is part of the i2cSlave opencores effort.
//// <http://www.opencores.org/cores//>                           ////
////                                                              ////
//// Module Description:                                          ////
//// You will need to modify this file to implement your 
//// interface.
//// Add your control and status bytes/bits to module inputs and outputs,
//// and also to the I2C read and write process blocks  
////                                                              ////
//// To Do:                                                       ////
//// 
////                                                              ////
//// Author(s):                                                   ////
//// - Steve Fielding, sfielding@base2designs.com                 ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
////                                                              ////
//// Copyright (C) 2008 Steve Fielding and OPENCORES.ORG          ////
////                                                              ////
//// This source file may be used and distributed without         ////
//// restriction provided that this copyright statement is not    ////
//// removed from the file and that any derivative work contains  ////
//// the original copyright notice and the associated disclaimer. ////
////                                                              ////
//// This source file is free software; you can redistribute it   ////
//// and/or modify it under the terms of the GNU Lesser General   ////
//// Public License as published by the Free Software Foundation; ////
//// either version 2.1 of the License, or (at your option) any   ////
//// later version.                                               ////
////                                                              ////
//// This source is distributed in the hope that it will be       ////
//// useful, but WITHOUT ANY WARRANTY; without even the implied   ////
//// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ////
//// PURPOSE. See the GNU Lesser General Public License for more  ////
//// details.                                                     ////
////                                                              ////
//// You should have received a copy of the GNU Lesser General    ////
//// Public License along with this source; if not, download it   ////
//// from <http://www.opencores.org/lgpl.shtml>                   ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
//
`include "i2cSlave_define.v"


module registerInterface (
  clk,
  addr,
  dataIn,
  writeEn,
  dataOut,
  reg0_auto_in,
  reg1_adc_cmd_out,
  reg2_ch0_upper_in,
  reg3_ch0_lower_in,
  reg4_ch1_upper_in,
  reg5_ch1_lower_in,
  reg6_ch2_upper_in,
  reg7_ch2_lower_in,
  reg8_ch3_upper_in,
  reg9_ch3_lower_in,
  reg10_ch4_upper_in,
  reg11_ch4_lower_in,
  reg12_ch5_upper_in,
  reg13_ch5_lower_in,
  //reg14_microphone_upper_in,
  //reg15_microphone_lower_in,
  //reg16_microphone_max_upper_in,
  //reg17_microphone_max_lower_in
);
input clk;
input [7:0] addr;
input [7:0] dataIn;
input writeEn;
output [7:0] dataOut;
input [7:0]  reg0_auto_in;
output [7:0] reg1_adc_cmd_out;
input [7:0]  reg2_ch0_upper_in;
input [7:0]  reg3_ch0_lower_in;
input [7:0]  reg4_ch1_upper_in;
input [7:0]  reg5_ch1_lower_in;
input [7:0]  reg6_ch2_upper_in;
input [7:0]  reg7_ch2_lower_in;
input [7:0]  reg8_ch3_upper_in;
input [7:0]  reg9_ch3_lower_in;
input [7:0]  reg10_ch4_upper_in;
input [7:0]  reg11_ch4_lower_in;
input [7:0]  reg12_ch5_upper_in;
input [7:0]  reg13_ch5_lower_in;
//input [7:0]  reg14_microphone_upper_in;
//input [7:0]  reg15_microphone_lower_in;
//input [7:0]  reg16_microphone_max_upper_in;
//input [7:0]  reg17_microphone_max_lower_in;

reg [7:0] dataOut;
reg [7:0] reg_auto;
reg [7:0] reg_adc_cmd;
reg [7:0] reg_ch0_upper;
reg [7:0] reg_ch0_lower;
reg [7:0] reg_ch1_upper;
reg [7:0] reg_ch1_lower;
reg [7:0] reg_ch2_upper;
reg [7:0] reg_ch2_lower;
reg [7:0] reg_ch3_upper;
reg [7:0] reg_ch3_lower;
reg [7:0] reg_ch4_upper;
reg [7:0] reg_ch4_lower;
reg [7:0] reg_ch5_upper;
reg [7:0] reg_ch5_lower;
//reg [7:0] reg_microphone_upper;
//reg [7:0] reg_microphone_lower;
//reg [7:0] reg_microphone_max_upper;
//reg [7:0] reg_microphone_max_lower;


// --- I2C Read
always @(posedge clk) begin
  case (addr)
    8'h00: dataOut <= reg_auto;  
    8'h01: dataOut <= reg_adc_cmd;
    8'h02: dataOut <= reg_ch0_upper;
    8'h03: dataOut <= reg_ch0_lower;
    8'h04: dataOut <= reg_ch1_upper;
    8'h05: dataOut <= reg_ch1_lower;
    8'h06: dataOut <= reg_ch2_upper;
    8'h07: dataOut <= reg_ch2_lower;
    8'h08: dataOut <= reg_ch3_upper;
    8'h09: dataOut <= reg_ch3_lower;
    8'h0a: dataOut <= reg_ch4_upper;
    8'h0b: dataOut <= reg_ch4_lower;
    8'h0c: dataOut <= reg_ch5_upper;
    8'h0d: dataOut <= reg_ch5_lower;
    //8'h0e: dataOut <= reg_microphone_upper;
    //8'h0f: dataOut <= reg_microphone_lower;
    //8'h10: dataOut <= reg_microphone_max_upper;
    //8'h11: dataOut <= reg_microphone_max_lower;
    default: dataOut <= 8'h00;
  endcase
end


// --- I2C Write (or update from GPIO state)
always @(posedge clk) begin

	//only reg_led writeable by I2C
  if (writeEn == 1'b1) begin
    case (addr)
      8'h01: reg_adc_cmd <= dataIn;
    endcase
  end
  	
  	//other regs update from GPIO state every clock
	reg_auto <= reg0_auto_in;
   reg_ch0_upper <= reg2_ch0_upper_in;
   reg_ch0_lower <= reg3_ch0_lower_in;
   reg_ch1_upper <= reg4_ch1_upper_in;
   reg_ch1_lower <= reg5_ch1_lower_in;
   reg_ch2_upper <= reg6_ch2_upper_in;
   reg_ch2_lower <= reg7_ch2_lower_in;
   reg_ch3_upper <= reg8_ch3_upper_in;
   reg_ch3_lower <= reg9_ch3_lower_in;
   reg_ch4_upper <= reg10_ch4_upper_in;
   reg_ch4_lower <= reg11_ch4_lower_in;
   reg_ch5_upper <= reg12_ch5_upper_in;
   reg_ch5_lower <= reg13_ch5_lower_in;
   //reg_microphone_upper <= reg14_microphone_upper_in;
   //reg_microphone_lower <= reg15_microphone_lower_in;
   //reg_microphone_max_upper <= reg16_microphone_max_upper_in;
   //reg_microphone_max_lower <= reg17_microphone_max_lower_in;
end

//assign reg1_led_out = reg_led;
assign reg1_adc_cmd_out = reg_adc_cmd;

endmodule


 
